1|W AH N
2|T UW
3|TH R IY
4|F AO R
4|F OW R
5|F AY V
6|S IH K S
7|S EH V AH N
8|EY T
9|N AY N
10|T EH N
11|IH L EH V AH N
12|T W EH L V
13|TH ER T IY N
14|F AO R T IY N
14|F OW R T IY N
15|F IH F T IY N
16|S IH K S T IY N
17|S EH V AH N T IY N
18|EY T IY N
19|N AY N T IY N
20|T W EH N T IY
30|TH ER D IY
40|F AO R T IY
40|F OW R T IY
50|F IH F T IY
60|S IH K S T IY
70|S EH V AH N T IY
80|EY T IY
90|N AY N T IY
100|W AH N HH AH N D R AH D
100|AH HH AH N D R AH D
hundred|HH AH N D R AH D
1000|W AH N TH AW Z AH N D
1000|AH TH AW Z AH N D
1,000|W AH N TH AW Z AH N D
1,000|AH TH AW Z AH N D
thousand|TH AW Z AH N D
1000000|W AH N M IH L Y AH N
1000000|AH M IH L Y AH N
1,000,000|W AH N M IH L Y AH N
1,000,000|AH M IH L Y AH N
million|M IH L Y AH N
and|AH N D
a|AH
